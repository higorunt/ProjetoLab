library verilog;
use verilog.vl_types.all;
entity ContadorCentesimosSegundo_vlg_vec_tst is
end ContadorCentesimosSegundo_vlg_vec_tst;
