library verilog;
use verilog.vl_types.all;
entity relogio_vlg_vec_tst is
end relogio_vlg_vec_tst;
