library verilog;
use verilog.vl_types.all;
entity ContadorSegundos_vlg_vec_tst is
end ContadorSegundos_vlg_vec_tst;
